module logic_xor (
    input logic a,
    input logic b,
    output logic y
);
    assign y = a ^ b; // Perform the XOR operation
endmodule
