module adder_32bit (input logic [31:0] a, b, output logic [31:0] z);

   assign z = a+b;

endmodule // sample
